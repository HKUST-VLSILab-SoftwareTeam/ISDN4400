`ifndef __SEVEN_SEG_DISPLAY_VH__
`define __SEVEN_SEG_DISPLAY_VH__

// 8'bABCDEFG(DP)
`define NUM_OFF     8'b11111111
`define NUM_0       8'b00000011
`define NUM_1       8'b10011111
`define NUM_2       8'b00100101
`define NUM_3       8'b00001101
`define NUM_4       8'b10011001
`define NUM_5       8'b01001001
`define NUM_6       8'b11000001
`define NUM_7       8'b00011111
`define NUM_8       8'b00000001
`define NUM_9       8'b00011001
`define NUM_A       8'b00010001
`define NUM_B       8'b11000001
`define NUM_C       8'b01100011
`define NUM_D       8'b10000101
`define NUM_E       8'b01100001
`define NUM_F       8'b00110001

`define AN0_ON      4'b1110
`define AN1_ON      4'b1101
`define AN2_ON      4'b1011
`define AN3_ON      4'b0111

`endif //__SEVEN_SEG_DISPLAY_H__

`ifndef __SEVEN_SEG_DISPLAY_VH__
`define __SEVEN_SEG_DISPLAY_VH__

`define NUM_OFF     8'b11111111
`define NUM_0       8'b00000011
`define NUM_1       8'b10011111
`define NUM_2       8'b10010010
`define NUM_3       8'b10000110
`define NUM_4       8'b11001100
`define NUM_5       8'b10100010
`define NUM_6       8'b11100000
`define NUM_7       8'b10001111
`define NUM_8       8'b10000000
`define NUM_9       8'b10001100
`define NUM_A       8'b10000100
`define NUM_B       8'b11100000
`define NUM_C       8'b10110001
`define NUM_D       8'b11000010
`define NUM_E       8'b10110000
`define NUM_F       8'b10011000

`define AN0_ON      4'b1110
`define AN1_ON      4'b1101
`define AN2_ON      4'b1011
`define AN3_ON      4'b0111

`endif //__SEVEN_SEG_DISPLAY_H__
